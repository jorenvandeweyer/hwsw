
module unsaved (
	clk_clk,
	resetn_reset_n,
	uart_0_external_rxd,
	uart_0_external_txd);	

	input		clk_clk;
	input		resetn_reset_n;
	input		uart_0_external_rxd;
	output		uart_0_external_txd;
endmodule
